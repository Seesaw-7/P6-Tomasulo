`ifndef __ISSUE_UNIT_SVH__
`define __ISSUE_UNIT_SVH__

`define ALU_LATE 1
`define BTU_LATE 1
`define MULT_LATE 9
`define LS_LATE 17

`endif 