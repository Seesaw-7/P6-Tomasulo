`ifndef __CACHE_SVH__
`define __CACHE_SVH__

`define CACHE_SIZE 256
`define CACHE_SIZE_BIT 8

`endif