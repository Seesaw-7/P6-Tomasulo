`ifndef __LS_UNIT_SVH__
`define __LS_UNIT_SVH__

`include "sys_defs.svh"
`include "dispatcher.svh"
`include "ls_queue.svh"

`endif
